--
--	The format of this file is proprietary information belonging
--	to Speed S.A. All copies of this file must include this notice.
--		Copyright (c) 1992,1993 and 1994 by SPEED S.A.
--

configuration SPDCH_AN2_CONF of SPDCH_AN2 is
	for SPDCH_AN2_ARCH
	end for;
end SPDCH_AN2_CONF;

configuration SPDCH_AN2_V_CONF of SPDCH_AN2_V is
	for SPDCH_AN2_V_ARCH
	end for;
end SPDCH_AN2_V_CONF;

configuration SPDCH_AN3_CONF of SPDCH_AN3 is
	for SPDCH_AN3_ARCH
	end for;
end SPDCH_AN3_CONF;

configuration SPDCH_AN3_V_CONF of SPDCH_AN3_V is
	for SPDCH_AN3_V_ARCH
	end for;
end SPDCH_AN3_V_CONF;

configuration SPDCH_AN4_CONF of SPDCH_AN4 is
	for SPDCH_AN4_ARCH
	end for;
end SPDCH_AN4_CONF;

configuration SPDCH_AN4_V_CONF of SPDCH_AN4_V is
	for SPDCH_AN4_V_ARCH
	end for;
end SPDCH_AN4_V_CONF;

configuration SPDCH_D12H_CONF of SPDCH_D12H is
	for SPDCH_D12H_ARCH
	end for;
end SPDCH_D12H_CONF;

configuration SPDCH_D24H_CONF of SPDCH_D24H is
	for SPDCH_D24H_ARCH
	end for;
end SPDCH_D24H_CONF;

configuration SPDCH_D38H_CONF of SPDCH_D38H is
	for SPDCH_D38H_ARCH
	end for;
end SPDCH_D38H_CONF;

configuration SPDCH_D12L_CONF of SPDCH_D12L is
	for SPDCH_D12L_ARCH
	end for;
end SPDCH_D12L_CONF;

configuration SPDCH_D24L_CONF of SPDCH_D24L is
	for SPDCH_D24L_ARCH
	end for;
end SPDCH_D24L_CONF;

configuration SPDCH_D38L_CONF of SPDCH_D38L is
	for SPDCH_D38L_ARCH
	end for;
end SPDCH_D38L_CONF;

configuration SPDCH_EN_CONF of SPDCH_EN is
	for SPDCH_EN_ARCH
	end for;
end SPDCH_EN_CONF;

configuration SPDCH_EN_V_CONF of SPDCH_EN_V is
	for SPDCH_EN_V_ARCH
	end for;
end SPDCH_EN_V_CONF;

configuration SPDCH_EO_CONF of SPDCH_EO is
	for SPDCH_EO_ARCH
	end for;
end SPDCH_EO_CONF;

configuration SPDCH_EO_V_CONF of SPDCH_EO_V is
	for SPDCH_EO_V_ARCH
	end for;
end SPDCH_EO_V_CONF;

configuration SPDCH_FA_CONF of SPDCH_FA is
	for SPDCH_FA_ARCH
	end for;
end SPDCH_FA_CONF;

configuration SPDCH_FD1_CONF of SPDCH_FD1 is
	for SPDCH_FD1_ARCH
	end for;
end SPDCH_FD1_CONF;

configuration SPDCH_FD2_CONF of SPDCH_FD2 is
	for SPDCH_FD2_ARCH
	end for;
end SPDCH_FD2_CONF;

configuration SPDCH_FD3_CONF of SPDCH_FD3 is
	for SPDCH_FD3_ARCH
	end for;
end SPDCH_FD3_CONF;

configuration SPDCH_FD4_CONF of SPDCH_FD4 is
        for SPDCH_FD4_ARCH
        end for;
end SPDCH_FD4_CONF;

configuration SPDCH_FD1_V_CONF of SPDCH_FD1_V is
	for SPDCH_FD1_V_ARCH
	end for;
end SPDCH_FD1_V_CONF;

configuration SPDCH_FD2_V_CONF of SPDCH_FD2_V is
	for SPDCH_FD2_V_ARCH
	end for;
end SPDCH_FD2_V_CONF;

configuration SPDCH_FD3_V_CONF of SPDCH_FD3_V is
	for SPDCH_FD3_V_ARCH
	end for;
end SPDCH_FD3_V_CONF;

configuration SPDCH_FD4_V_CONF of SPDCH_FD4_V is
        for SPDCH_FD4_V_ARCH
        end for;
end SPDCH_FD4_V_CONF;

configuration SPDCH_FJK1_CONF of SPDCH_FJK1 is
	for SPDCH_FJK1_ARCH
	end for;
end SPDCH_FJK1_CONF;

configuration SPDCH_FJK2_CONF of SPDCH_FJK2 is
	for SPDCH_FJK2_ARCH
	end for;
end SPDCH_FJK2_CONF;

configuration SPDCH_FJK3_CONF of SPDCH_FJK3 is
	for SPDCH_FJK3_ARCH
	end for;
end SPDCH_FJK3_CONF;

configuration SPDCH_FJK4_CONF of SPDCH_FJK4 is
        for SPDCH_FJK4_ARCH
        end for;
end SPDCH_FJK4_CONF;

configuration SPDCH_GND_CONF of SPDCH_GND is
	for SPDCH_GND_ARCH
	end for;
end SPDCH_GND_CONF;

configuration SPDCH_GND_V_CONF of SPDCH_GND_V is
	for SPDCH_GND_V_ARCH
	end for;
end SPDCH_GND_V_CONF;

configuration SPDCH_HA_CONF of SPDCH_HA is
	for SPDCH_HA_ARCH
	end for;
end SPDCH_HA_CONF;

configuration SPDCH_IV_CONF of SPDCH_IV is
	for SPDCH_IV_ARCH
	end for;
end SPDCH_IV_CONF;

configuration SPDCH_IV_V_CONF of SPDCH_IV_V is
	for SPDCH_IV_V_ARCH
	end for;
end SPDCH_IV_V_CONF;

configuration SPDCH_LD1_CONF of SPDCH_LD1 is
	for SPDCH_LD1_ARCH
	end for;
end SPDCH_LD1_CONF;

configuration SPDCH_LD2_CONF of SPDCH_LD2 is
	for SPDCH_LD2_ARCH
	end for;
end SPDCH_LD2_CONF;

configuration SPDCH_LD3_CONF of SPDCH_LD3 is
	for SPDCH_LD3_ARCH
	end for;
end SPDCH_LD3_CONF;

configuration SPDCH_LD4_CONF of SPDCH_LD4 is
	for SPDCH_LD4_ARCH
	end for;
end SPDCH_LD4_CONF;

configuration SPDCH_LD5_CONF of SPDCH_LD5 is
	for SPDCH_LD5_ARCH
	end for;
end SPDCH_LD5_CONF;

configuration SPDCH_LD6_CONF of SPDCH_LD6 is
	for SPDCH_LD6_ARCH
	end for;
end SPDCH_LD6_CONF;

configuration SPDCH_LD7_CONF of SPDCH_LD7 is
	for SPDCH_LD7_ARCH
	end for;
end SPDCH_LD7_CONF;

configuration SPDCH_LD8_CONF of SPDCH_LD8 is
	for SPDCH_LD8_ARCH
	end for;
end SPDCH_LD8_CONF;

configuration SPDCH_LD1_V_CONF of SPDCH_LD1_V is
	for SPDCH_LD1_V_ARCH
	end for;
end SPDCH_LD1_V_CONF;

configuration SPDCH_LD2_V_CONF of SPDCH_LD2_V is
	for SPDCH_LD2_V_ARCH
	end for;
end SPDCH_LD2_V_CONF;

configuration SPDCH_LD3_V_CONF of SPDCH_LD3_V is
	for SPDCH_LD3_V_ARCH
	end for;
end SPDCH_LD3_V_CONF;

configuration SPDCH_LD4_V_CONF of SPDCH_LD4_V is
	for SPDCH_LD4_V_ARCH
	end for;
end SPDCH_LD4_V_CONF;

configuration SPDCH_LD5_V_CONF of SPDCH_LD5_V is
	for SPDCH_LD5_V_ARCH
	end for;
end SPDCH_LD5_V_CONF;

configuration SPDCH_LD6_V_CONF of SPDCH_LD6_V is
	for SPDCH_LD6_V_ARCH
	end for;
end SPDCH_LD6_V_CONF;

configuration SPDCH_LD7_V_CONF of SPDCH_LD7_V is
	for SPDCH_LD7_V_ARCH
	end for;
end SPDCH_LD7_V_CONF;

configuration SPDCH_LD8_V_CONF of SPDCH_LD8_V is
	for SPDCH_LD8_V_ARCH
	end for;
end SPDCH_LD8_V_CONF;

configuration SPDCH_LSRA_CONF of SPDCH_LSRA is
	for SPDCH_LSRA_ARCH
	end for;
end SPDCH_LSRA_CONF;

configuration SPDCH_LSRB_CONF of SPDCH_LSRB is
	for SPDCH_LSRB_ARCH
	end for;
end SPDCH_LSRB_CONF;

configuration SPDCH_MX21_CONF of SPDCH_MX21 is
	for SPDCH_MX21_ARCH
	end for;
end SPDCH_MX21_CONF;

configuration SPDCH_MX21_V_CONF of SPDCH_MX21_V is
	for SPDCH_MX21_V_ARCH
	end for;
end SPDCH_MX21_V_CONF;

configuration SPDCH_MX41_CONF of SPDCH_MX41 is
	for SPDCH_MX41_ARCH
	end for;
end SPDCH_MX41_CONF;

configuration SPDCH_MX41_V_CONF of SPDCH_MX41_V is
	for SPDCH_MX41_V_ARCH
	end for;
end SPDCH_MX41_V_CONF;

configuration SPDCH_ND2_CONF of SPDCH_ND2 is
	for SPDCH_ND2_ARCH
	end for;
end SPDCH_ND2_CONF;

configuration SPDCH_ND2_V_CONF of SPDCH_ND2_V is
	for SPDCH_ND2_V_ARCH
	end for;
end SPDCH_ND2_V_CONF;

configuration SPDCH_ND3_CONF of SPDCH_ND3 is
	for SPDCH_ND3_ARCH
	end for;
end SPDCH_ND3_CONF;

configuration SPDCH_ND3_V_CONF of SPDCH_ND3_V is
	for SPDCH_ND3_V_ARCH
	end for;
end SPDCH_ND3_V_CONF;

configuration SPDCH_ND4_CONF of SPDCH_ND4 is
	for SPDCH_ND4_ARCH
	end for;
end SPDCH_ND4_CONF;

configuration SPDCH_ND4_V_CONF of SPDCH_ND4_V is
	for SPDCH_ND4_V_ARCH
	end for;
end SPDCH_ND4_V_CONF;

configuration SPDCH_NOP_CONF of SPDCH_NOP is
	for SPDCH_NOP_ARCH
	end for;
end SPDCH_NOP_CONF;

configuration SPDCH_NOP_V_CONF of SPDCH_NOP_V is
	for SPDCH_NOP_V_ARCH
	end for;
end SPDCH_NOP_V_CONF;

configuration SPDCH_NR2_CONF of SPDCH_NR2 is
	for SPDCH_NR2_ARCH
	end for;
end SPDCH_NR2_CONF;

configuration SPDCH_NR2_V_CONF of SPDCH_NR2_V is
	for SPDCH_NR2_V_ARCH
	end for;
end SPDCH_NR2_V_CONF;

configuration SPDCH_NR3_CONF of SPDCH_NR3 is
	for SPDCH_NR3_ARCH
	end for;
end SPDCH_NR3_CONF;

configuration SPDCH_NR3_V_CONF of SPDCH_NR3_V is
	for SPDCH_NR3_V_ARCH
	end for;
end SPDCH_NR3_V_CONF;

configuration SPDCH_NR4_CONF of SPDCH_NR4 is
	for SPDCH_NR4_ARCH
	end for;
end SPDCH_NR4_CONF;

configuration SPDCH_NR4_V_CONF of SPDCH_NR4_V is
	for SPDCH_NR4_V_ARCH
	end for;
end SPDCH_NR4_V_CONF;

configuration SPDCH_OR2_CONF of SPDCH_OR2 is
	for SPDCH_OR2_ARCH
	end for;
end SPDCH_OR2_CONF;

configuration SPDCH_OR2_V_CONF of SPDCH_OR2_V is
	for SPDCH_OR2_V_ARCH
	end for;
end SPDCH_OR2_V_CONF;

configuration SPDCH_OR3_CONF of SPDCH_OR3 is
	for SPDCH_OR3_ARCH
	end for;
end SPDCH_OR3_CONF;

configuration SPDCH_OR3_V_CONF of SPDCH_OR3_V is
	for SPDCH_OR3_V_ARCH
	end for;
end SPDCH_OR3_V_CONF;

configuration SPDCH_OR4_CONF of SPDCH_OR4 is
	for SPDCH_OR4_ARCH
	end for;
end SPDCH_OR4_CONF;

configuration SPDCH_OR4_V_CONF of SPDCH_OR4_V is
	for SPDCH_OR4_V_ARCH
	end for;
end SPDCH_OR4_V_CONF;

configuration SPDCH_PD_CONF of SPDCH_PD is
	for SPDCH_PD_ARCH
	end for;
end SPDCH_PD_CONF;

configuration SPDCH_PU_CONF of SPDCH_PU is
	for SPDCH_PU_ARCH
	end for;
end SPDCH_PU_CONF;

configuration SPDCH_VDD_CONF of SPDCH_VDD is
	for SPDCH_VDD_ARCH
	end for;
end SPDCH_VDD_CONF;

configuration SPDCH_VDD_V_CONF of SPDCH_VDD_V is
	for SPDCH_VDD_V_ARCH
	end for;
end SPDCH_VDD_V_CONF;
