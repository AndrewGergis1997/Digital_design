//---------------------------------------------------------------------------
// svassist_pkg
//
//   A package that contains the functions needed to generate
//   the dynamic hierarchy and connectivity of a UVM environment.
//
//   Version: 3.0 - Re-written for UVM 1.0 use only. 
//                  No changes required to UVM library 
//
//
//   Copyright Mentor Graphics Corporation, 2007-2011. 
//   All Rights Reserved.
//   UNPUBLISHED, LICENSED SOFTWARE. CONFIDENTIAL AND PROPRIETARY INFORMATION
//   WHICH IS THE PROPERTY OF MENTOR GRAPHICS CORPORATION OR ITS LICENSORS.
//---------------------------------------------------------------------------

`ifndef SVASSIST_PKG_SV
`define SVASSIST_PKG_SV

package svassist_pkg;
import uvm_pkg::*;

  `include "svassist_inc.svp"

endpackage: svassist_pkg

`endif