-- Copyright Mentor Graphics Corporation 2004
--
--    All Rights Reserved.
--
-- THIS WORK CONTAINS TRADE SECRET
-- AND PROPRIETARY INFORMATION WHICH IS THE
-- PROPERTY OF MENTOR GRAPHICS
-- CORPORATION OR ITS LICENSORS AND IS
-- SUBJECT TO LICENSE TERMS. 

--**************************************************************************
--**
--**
--**************************************************************************
--- *************************************************************************

library ieee;
use     ieee.std_logic_1164.all;
use 	IEEE.std_logic_arith.all;

library work;
use 	work.amba.all;
-- use 	work.ahb_iface_pkg.all ;
-- use 	work.bbcreg_pkg.all ;
-- use 	work.bbc_sram_pkg.all ;
-- use 	work.bbc_intc_pkg.all ;
--!!!!!!!!!!!!!!!!!!!!!!!!!!!! begin of BBCDesigned generated part !!!!!!!!!!!!
-- import generated packages for bus interfaces
--$BBCDesigner: BIF packages$
--!!!!!!!!!!!!!!!!!!!!!!!!!!!! end of BBCDesigned generated part !!!!!!!!!!!!

-------------------------------------------------------------------------------
--  entity of bbc_top  declaration
-------------------------------------------------------------------------------
entity bbc_top is

  port (
  
--!!!!!!!!!!!!!!!!!!!!!!!!!!!! begin of BBCDesigned generated part !!!!!!!!!!!!
--$BBCDesigner: top signals list$
--!!!!!!!!!!!!!!!!!!!!!!!!!!!! end of BBCDesigned generated part !!!!!!!!!!!!

--    DUMMYDUMMYDUMMY  :   in Std_Logic                         -- dummy signal
    );

end bbc_top ;


architecture structural of bbc_top is

begin

--!!!!!!!!!!!!!!!!!!!!!!!!!!!! begin of BBCDesigned generated part !!!!!!!!!!!!
--$BBCDesigner: top components list$
--!!!!!!!!!!!!!!!!!!!!!!!!!!!! end of BBCDesigned generated part !!!!!!!!!!!!

end structural ;




