//------------------------------------------------------------------------------
//   Copyright 2010 Mentor Graphics Corporation
//
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------------------------
class ready_valid_sequence_item extends ovm_sequence_item;
  `ovm_object_utils( ready_valid_sequence_item );

  bit [7:0] m_data;

  function new( string name = "" );
    super.new( name );
  endfunction

  function void do_print( ovm_printer printer );
    printer.print_string("Type" , "Ready Valid Transaction" );
    printer.print_field("Data" , m_data , $bits( m_data ) );
  endfunction

  function bit do_compare( ovm_object rhs , ovm_comparer comparer );
    ready_valid_sequence_item t;

    assert( $cast( t , rhs ) );
    return m_data == t.m_data;
  endfunction

endclass
