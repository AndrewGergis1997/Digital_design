// $Id: //dvt/vtech/dev/6.4x/avm/libraries/systemverilog/avm/utils/code/avm_utils.svh#3 $
//----------------------------------------------------------------------
//   Copyright 2005-2008 Mentor Graphics Corporation
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------

`include "utils/avm_threaded_component.svh"
`include "utils/avm_env.svh"

`include "utils/avm_pair.svh"
`include "utils/avm_in_order_comparator.svh"
`include "utils/avm_algorithmic_comparator.svh"

`include "utils/avm_random_stimulus.svh"
`include "utils/avm_subscriber.svh"


